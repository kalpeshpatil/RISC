library verilog;
use verilog.vl_types.all;
entity controller is
    generic(
        fetch1          : integer := 0;
        fetch2          : integer := 1;
        fetch_check     : integer := 2;
        add1            : integer := 3;
        add2            : integer := 4;
        add3            : integer := 5;
        adi1            : integer := 7;
        adi2            : integer := 8;
        adi3            : integer := 9;
        nan             : integer := 6;
        lhi1            : integer := 10;
        lhi2            : integer := 11;
        sl1             : integer := 12;
        sl2             : integer := 13;
        sl3             : integer := 14;
        sl4             : integer := 15;
        sl5             : integer := 16;
        sl6             : integer := 17;
        slm             : integer := 18;
        l1              : integer := 19;
        l2              : integer := 20;
        l3              : integer := 21;
        s1              : integer := 22;
        s2              : integer := 23;
        s3              : integer := 24;
        beq1            : integer := 25;
        beq2            : integer := 26;
        beq3            : integer := 27;
        beq4            : integer := 28;
        jalr            : integer := 29;
        jal1            : integer := 30;
        jal2            : integer := 31;
        jlr1            : integer := 32;
        jlr2            : integer := 33;
        jump            : integer := 34;
        updater         : integer := 35;
        beqcheck        : integer := 36
    );
    port(
        clock           : in     vl_logic;
        clock_50        : in     vl_logic;
        curr_state      : out    vl_logic_vector(5 downto 0);
        reg_7           : out    vl_logic_vector(15 downto 0);
        reg_6           : out    vl_logic_vector(15 downto 0);
        edb_out         : out    vl_logic_vector(15 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of fetch1 : constant is 1;
    attribute mti_svvh_generic_type of fetch2 : constant is 1;
    attribute mti_svvh_generic_type of fetch_check : constant is 1;
    attribute mti_svvh_generic_type of add1 : constant is 1;
    attribute mti_svvh_generic_type of add2 : constant is 1;
    attribute mti_svvh_generic_type of add3 : constant is 1;
    attribute mti_svvh_generic_type of adi1 : constant is 1;
    attribute mti_svvh_generic_type of adi2 : constant is 1;
    attribute mti_svvh_generic_type of adi3 : constant is 1;
    attribute mti_svvh_generic_type of nan : constant is 1;
    attribute mti_svvh_generic_type of lhi1 : constant is 1;
    attribute mti_svvh_generic_type of lhi2 : constant is 1;
    attribute mti_svvh_generic_type of sl1 : constant is 1;
    attribute mti_svvh_generic_type of sl2 : constant is 1;
    attribute mti_svvh_generic_type of sl3 : constant is 1;
    attribute mti_svvh_generic_type of sl4 : constant is 1;
    attribute mti_svvh_generic_type of sl5 : constant is 1;
    attribute mti_svvh_generic_type of sl6 : constant is 1;
    attribute mti_svvh_generic_type of slm : constant is 1;
    attribute mti_svvh_generic_type of l1 : constant is 1;
    attribute mti_svvh_generic_type of l2 : constant is 1;
    attribute mti_svvh_generic_type of l3 : constant is 1;
    attribute mti_svvh_generic_type of s1 : constant is 1;
    attribute mti_svvh_generic_type of s2 : constant is 1;
    attribute mti_svvh_generic_type of s3 : constant is 1;
    attribute mti_svvh_generic_type of beq1 : constant is 1;
    attribute mti_svvh_generic_type of beq2 : constant is 1;
    attribute mti_svvh_generic_type of beq3 : constant is 1;
    attribute mti_svvh_generic_type of beq4 : constant is 1;
    attribute mti_svvh_generic_type of jalr : constant is 1;
    attribute mti_svvh_generic_type of jal1 : constant is 1;
    attribute mti_svvh_generic_type of jal2 : constant is 1;
    attribute mti_svvh_generic_type of jlr1 : constant is 1;
    attribute mti_svvh_generic_type of jlr2 : constant is 1;
    attribute mti_svvh_generic_type of jump : constant is 1;
    attribute mti_svvh_generic_type of updater : constant is 1;
    attribute mti_svvh_generic_type of beqcheck : constant is 1;
end controller;
