library verilog;
use verilog.vl_types.all;
entity se6_16 is
    port(
        \in\            : in     vl_logic_vector(5 downto 0);
        \out\           : out    vl_logic_vector(15 downto 0)
    );
end se6_16;
